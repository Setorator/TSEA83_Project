-----------------------------------------
------------BLOCK_RAM--------------------
-----------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;                        -- IEEE library for the unsigned type
                                                 -- and various arithmetic operations


entity RAM is
	port (
		clk			: in std_logic;					-- Clock pulse
		
		-- port 1
		x1 			: in unsigned(5 downto 0);					-- 64 columns, only 40 is used
		y1 			: in unsigned(4 downto 0);					-- 32 rows, only 30 used
		we 			: in std_logic;								-- Write enable
		data1			: in std_logic_vector(1 downto 0);		-- Data to be written (tile-type)

		-- port 2
		x2 			: in unsigned(5 downto 0);					-- 64 columns, only 40 is used
		y2 			: in unsigned(4 downto 0);					-- 32 rows, only 30 used
		re 			: in std_logic;								-- Read enable
		data2			: out std_logic_vector(1 downto 0)		-- Data to be read (tile-type)
	);
end RAM;

architecture Behavioral of RAM is

	-- Declaration of a two-port RAM
	-- with 2048 adresses and 8 bits width
	-- (We only uses 40*30 = 1200 adresses,
	-- each containing a 8-bit colour.)
	type ram_t is array(0 to 2047) of 
		std_logic_vector(1 downto 0);
	
	-- Set all bits to zero
	signal ram : ram_t := ( "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00", others => (others => '1'));
	
	begin
	
	
	process(clk)
	begin
		if rising_edge(clk) then
		
			-- Synched write port 1
			if (we = '0') then
				ram(30*to_integer(y1)+
					to_integer(x1)) <= data1;
			end if;
		
			-- synched read from port 2
			if (re = '0') then 
				data2 <= ram(30*to_integer(y2)+
									to_integer(x2));
			end if;
		
		end if;
	end process;
	
end Behavioral;
	
	
	
