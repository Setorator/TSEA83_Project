-----------------------------------------
------------BLOCK_RAM--------------------
-----------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;                        -- IEEE library for the unsigned type
                                                 -- and various arithmetic operations


entity RAM is
	port (
		clk			: in std_logic;					-- Clock pulse
		rst			: in std_logic;					-- Reset 						-- Never used???
		
		-- port 1 (write)
		x_write 		: in unsigned(5 downto 0);					-- 64 columns, only 40 is used
		y_write		: in unsigned(4 downto 0);					-- 32 rows, only 30 used
		we 			: in std_logic;								-- Write enable
		data_write	: in std_logic_vector(1 downto 0);		-- Data to be written (tile-type)

		-- port 2 (read)
		x_read		: in unsigned(5 downto 0);					-- 64 columns, only 40 is used
		y_read		: in unsigned(4 downto 0);					-- 32 rows, only 30 used
		re 			: in std_logic;								-- Read enable
		data_read	: out std_logic_vector(1 downto 0)		-- Data to be read (tile-type)
		
	);
end RAM;

architecture Behavioral of RAM is


	-- Declaration of a two-port RAM
	-- with 1200 adresses, each containing a 2-bit tile_type.
	type ram_t is array(0 to 1199) of 
		std_logic_vector(1 downto 0);
		
-- 	The ram only contains a 2-bit binary-code of the specific tile type on 
-- 	the corresponding position. The color is later given in the PIX_GEN module
--		This is to minimize the space required, since 2 bits (tile type) < 8 bits (color)


	-- ("00", "01", "10", "11") = (Floor, Food, Undefined, Wall)
	signal ram : ram_t := ( "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00", 
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									
									"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
									"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11", 
									"11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01", 
									"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","11", -- Row 8
									"11","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11", 
									"11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","11", 
									"11","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11","11","00",
									
									"00","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","00",
									
									"00","11","11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","01", 
									"01","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11","11","00",
									
									"11","11","11","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","00", 
									"00","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","11","11","11",
									
									"00","00","01","01","01","01","01","01","01","01","01","01","01","11","00","00","00","00","00","00", 
									"00","00","00","00","00","00","11","01","01","01","01","01","01","01","01","01","01","01","00","00",
									
									"11","11","11","11","11","11","11","11","11","01","11","11","01","11","00","00","00","00","00","00", 
									"00","00","00","00","00","00","11","01","11","11","01","11","11","11","11","11","11","11","11","11",
									
									"00","11","11","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","11", -- Row 16
									"11","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","11","11","00",
									
									"00","11","11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","01", 
									"01","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11", 
									"11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","01","01","01","01","01","01","01","01","01","11", 
									"11","01","01","01","01","01","01","01","01","01","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","01","01","01","01","11","11","01","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","01","11","11","01","01","01","01","01","11","00",
									
									"00","11","11","11","11","11","01","11","11","01","01","01","01","01","01","01","01","01","01","01", 
									"01","01","01","01","01","01","01","01","01","01","01","11","11","01","11","11","11","11","11","00",
									
									"00","11","11","11","11","11","01","11","11","01","11","11","11","11","11","11","11","11","11","11", 
									"11","11","11","11","11","11","11","11","11","11","01","11","11","01","11","11","11","11","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11", -- Row 24
									"11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","01","11", 
									"11","01","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","01","11","00",
									
									"00","11","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01", 
									"01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","11","00",
									
									"00","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11",
									"11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","11","00",
									
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00", 
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
									
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00", 
									"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00", others => (others => '0'));
									
	
	begin


	
	-- Our read and write process for the ram.
	Read_Write : process(clk)
	begin
		if rising_edge(clk) then	
			if (rst = '0') then
				-- Synched write port 1	
				if (we = '0') then
					ram(40*to_integer(y_write) + to_integer(x_write)) <= data_write;
				end if;
		
				-- synched read from port 2
				if (re = '0') then 
					data_read <= ram(40*to_integer(y_read) + to_integer(x_read));
				end if;
			end if;
		end if;
	end process;
	
end Behavioral;
	
	
	
